LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TEST_BENCH IS 
END ENTITY;

ARCHITECTURE TB OF TEST_BENCH IS
SIGNAL S: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL F: STD_LOGIC_VECTOR(250 DOWNTO 0);
BEGIN
UUT: ENTITY WORK.DECODER_8IP PORT MAP(S,F);
S<="00000000","11111111" AFTER 300 NS,"11010111" AFTER 600 NS,"10101010" AFTER 900 NS,"01001011" AFTER 2000 NS;
END ARCHITECTURE;