LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODER_8IP IS
GENERIC(
I: NATURAL := 8;
O: NATURAL := 251
);
PORT(
A: IN STD_LOGIC_VECTOR(I-1 DOWNTO 0);
F: OUT STD_LOGIC_VECTOR(O-1 DOWNTO 0)
);
END ENTITY;


ARCHITECTURE STRUC OF DECODER_8IP IS
SIGNAL S: STD_LOGIC_VECTOR(I-1 DOWNTO 0);

--COMPONENT DECLARATION
COMPONENT AND_8IP
GENERIC(
n: NATURAL:=8
);
PORT(
A: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
F: OUT STD_LOGIC
);
END COMPONENT;

-- BEGINIGN SEQUENTIAL SENTENCES
BEGIN
PROCESS(A)
VARIABLE VAR:INTEGER:=0;
BEGIN
FOR VAR IN (I-1) DOWNTO 0 LOOP
S(VAR)<=(NOT A(VAR));
END LOOP;
END PROCESS;
AND0: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(0));
AND1: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(1));
AND2: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(2));
AND3: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(3));
AND4: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(4));
AND5: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(5));
AND6: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(6));
AND7: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(7));
AND8: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(8));
AND9: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(9));
AND10: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(10));
AND11: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(11));
AND12: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(12));
AND13: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(13));
AND14: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(14));
AND15: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(15));
AND16: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(16));
AND17: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(17));
AND18: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(18));
AND19: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(19));
AND20: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(20));
AND21: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(21));
AND22: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(22));
AND23: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(23));
AND24: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(24));
AND25: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(25));
AND26: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(26));
AND27: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(27));
AND28: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(28));
AND29: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(29));
AND30: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(30));
AND31: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(31));
AND32: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(32));
AND33: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(33));
AND34: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(34));
AND35: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(35));
AND36: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(36));
AND37: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(37));
AND38: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(38));
AND39: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(39));
AND40: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(40));
AND41: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(41));
AND42: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(42));
AND43: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(43));
AND44: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(44));
AND45: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(45));
AND46: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(46));
AND47: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(47));
AND48: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(48));
AND49: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(49));
AND50: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(50));
AND51: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(51));
AND52: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(52));
AND53: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(53));
AND54: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(54));
AND55: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(55));
AND56: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(56));
AND57: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(57));
AND58: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(58));
AND59: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(59));
AND60: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(60));
AND61: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(61));
AND62: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(62));
AND63: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(63));
AND64: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(64));
AND65: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(65));
AND66: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(66));
AND67: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(67));
AND68: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(68));
AND69: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(69));
AND70: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(70));
AND71: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(71));
AND72: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(72));
AND73: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(73));
AND74: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(74));
AND75: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(75));
AND76: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(76));
AND77: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(77));
AND78: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(78));
AND79: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(79));
AND80: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(80));
AND81: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(81));
AND82: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(82));
AND83: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(83));
AND84: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(84));
AND85: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(85));
AND86: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(86));
AND87: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(87));
AND88: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(88));
AND89: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(89));
AND90: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(90));
AND91: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(91));
AND92: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(92));
AND93: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(93));
AND94: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(94));
AND95: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(95));
AND96: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(96));
AND97: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(97));
AND98: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(98));
AND99: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(99));
AND100: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(100));
AND101: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(101));
AND102: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(102));
AND103: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(103));
AND104: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(104));
AND105: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(105));
AND106: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(106));
AND107: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(107));
AND108: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(108));
AND109: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(109));
AND110: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(110));
AND111: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(111));
AND112: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(112));
AND113: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(113));
AND114: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(114));
AND115: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(115));
AND116: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(116));
AND117: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(117));
AND118: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(118));
AND119: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(119));
AND120: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(120));
AND121: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(121));
AND122: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(122));
AND123: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(123));
AND124: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(124));
AND125: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(125));
AND126: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(126));
AND127: AND_8IP PORT MAP(A(7)=>S(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(127));
AND128: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(128));
AND129: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(129));
AND130: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(130));
AND131: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(131));
AND132: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(132));
AND133: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(133));
AND134: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(134));
AND135: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(135));
AND136: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(136));
AND137: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(137));
AND138: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(138));
AND139: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(139));
AND140: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(140));
AND141: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(141));
AND142: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(142));
AND143: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(143));
AND144: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(144));
AND145: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(145));
AND146: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(146));
AND147: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(147));
AND148: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(148));
AND149: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(149));
AND150: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(150));
AND151: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(151));
AND152: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(152));
AND153: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(153));
AND154: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(154));
AND155: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(155));
AND156: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(156));
AND157: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(157));
AND158: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(158));
AND159: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(159));
AND160: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(160));
AND161: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(161));
AND162: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(162));
AND163: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(163));
AND164: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(164));
AND165: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(165));
AND166: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(166));
AND167: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(167));
AND168: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(168));
AND169: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(169));
AND170: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(170));
AND171: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(171));
AND172: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(172));
AND173: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(173));
AND174: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(174));
AND175: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(175));
AND176: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(176));
AND177: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(177));
AND178: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(178));
AND179: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(179));
AND180: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(180));
AND181: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(181));
AND182: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(182));
AND183: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(183));
AND184: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(184));
AND185: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(185));
AND186: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(186));
AND187: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(187));
AND188: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(188));
AND189: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(189));
AND190: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(190));
AND191: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>S(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(191));
AND192: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(192));
AND193: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(193));
AND194: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(194));
AND195: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(195));
AND196: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(196));
AND197: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(197));
AND198: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(198));
AND199: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(199));
AND200: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(200));
AND201: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(201));
AND202: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(202));
AND203: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(203));
AND204: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(204));
AND205: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(205));
AND206: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(206));
AND207: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(207));
AND208: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(208));
AND209: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(209));
AND210: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(210));
AND211: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(211));
AND212: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(212));
AND213: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(213));
AND214: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(214));
AND215: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(215));
AND216: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(216));
AND217: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(217));
AND218: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(218));
AND219: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(219));
AND220: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(220));
AND221: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(221));
AND222: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(222));
AND223: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>S(5),A(4)=>A(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(223));
AND224: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(224));
AND225: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(225));
AND226: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(226));
AND227: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(227));
AND228: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(228));
AND229: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(229));
AND230: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(230));
AND231: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(231));
AND232: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(232));
AND233: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(233));
AND234: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(234));
AND235: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(235));
AND236: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(236));
AND237: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(237));
AND238: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(238));
AND239: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>S(4),A(3)=>A(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(239));
AND240: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(240));
AND241: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(241));
AND242: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(242));
AND243: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>S(2),A(1)=>A(1),A(0)=>A(0),F=>F(243));
AND244: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>S(0),F=>F(244));
AND245: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>S(1),A(0)=>A(0),F=>F(245));
AND246: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>S(0),F=>F(246));
AND247: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>S(3),A(2)=>A(2),A(1)=>A(1),A(0)=>A(0),F=>F(247));
AND248: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>S(0),F=>F(248));
AND249: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>S(1),A(0)=>A(0),F=>F(249));
AND250: AND_8IP PORT MAP(A(7)=>A(7),A(6)=>A(6),A(5)=>A(5),A(4)=>A(4),A(3)=>A(3),A(2)=>S(2),A(1)=>A(1),A(0)=>S(0),F=>F(250));
END ARCHITECTURE;




