LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TEST_BENCH IS 
END ENTITY;

ARCHITECTURE TB OF TEST_BENCH IS
SIGNAL S: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL F: STD_LOGIC;
BEGIN
UUT: ENTITY WORK.AND_8IP PORT MAP(A=>S,F=>F);
S<="11110011","00000000" AFTER 10 NS,"11111111" AFTER 20NS,"01010101" AFTER 50 NS;
END ARCHITECTURE;