LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AND_8IP IS
GENERIC(
n: NATURAL:=8
);
PORT(
A: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0):="00000000";
F: OUT STD_LOGIC
);
END ENTITY;

ARCHITECTURE DF OF AND_8IP IS
BEGIN
F<=(A(0) AND A(1) AND A(2) AND A(3) AND A(4) AND A(5) AND A(6) AND A(7));
END ARCHITECTURE;
